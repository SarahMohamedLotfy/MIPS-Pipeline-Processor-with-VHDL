library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity Instrcontroller is
port(
    tag :in std_logic_vector(2 downto 0);
    index : in std_logic_vector(4 downto 0); -- to select which group.
    clk,rst,rd,memory_ready : in std_logic;-- ready signal from main memory to indicate that transfering data between main memory and cache is done

    Cache_read,Cache_Bus_Write,Memory_Bus_Read,Cache_Bus_Read,Memory_Bus_Write: out std_logic;
    hit_miss,Stall :out std_logic --Hit =1 miss =0
);
end Instrcontroller;


architecture controller_arch of Instrcontroller is


type states is (start, read_Hit,read_miss,Write_Back,Read_Main);
signal current_state : states := start;

    signal ReadMissSignal:std_logic; --to indicate that the state read main is coming from read miss
    signal sig_wr : std_logic;
    signal sig_rd : std_logic;
    signal sig_dbin : std_logic;
    signal sig_vdin : std_logic;
    signal sig_tagin : std_logic_vector(2 downto 0);
    signal sig_dbout : std_logic;
    signal sig_vdout : std_logic;
    signal sig_tagout : std_logic_vector(2 downto 0);
    
    begin
    
        f0:entity work.TVD port map(index, clk ,sig_wr ,sig_rd ,sig_tagin ,sig_dbin ,sig_vdin ,sig_tagout ,sig_dbout ,sig_vdout);

--Decide state process
DecideState : process(clk,rst)
begin
      if rst = '1' then
            current_state <= start;
      elsif rising_edge(clk) then 
        case current_state is
            when start =>
                if(rd = '1' )then----------------->>>>>>>>Read
                    if(tag = sig_tagout and sig_vdout = '1')then----------------->>>>>>>>> Hit
                    current_state <= read_Hit; 
                    else------------>>>>> Miss
                    current_state <= read_miss;
                    end if;
                end if;
            when read_miss =>
                if (sig_vdout = '1' and sig_dbout='1' ) then current_state <= Write_Back; else current_state <=Read_Main ; end if;
            
            when read_Hit=>
                current_state<=start;
            when Read_Main =>
                if memory_ready='1' and ReadMissSignal ='1'  then
                    current_state <= read_Hit;
                end if;
            when  Write_Back=>
                if memory_ready='1' then current_state <= Read_Main ;end if;
        end case;
      end if;
end process ; -- DecideState
StatesOutput:process (current_state,rd,tag,sig_tagout,sig_vdout,memory_ready) 
begin
    case current_state is
        when start =>
        ReadMissSignal <='0';
        sig_tagin<=tag; 
        sig_wr<='0' ;sig_rd<='1';
        Cache_read<='0';Cache_Bus_Write<='0';Memory_Bus_Read<='0';Cache_Bus_Read<='0';Memory_Bus_Write<='0';
        hit_miss<='0';Stall<='0';

        when read_Hit =>
        ReadMissSignal <='0';
        sig_tagin<=tag;
        sig_wr<='0' ;sig_rd<='0';
        Cache_read<='1'; Cache_Bus_Write<='0';Memory_Bus_Read<='0';Cache_Bus_Read<='0';Memory_Bus_Write<='0';
        hit_miss<='1';Stall<='0';

        when read_miss =>
        ReadMissSignal <='1';
        sig_tagin<=tag;
        sig_wr<='0' ;sig_rd<='0';
      
        Cache_read<='0'; Cache_Bus_Write<='0';Memory_Bus_Read<='0';Cache_Bus_Read<='0';Memory_Bus_Write<='0';
        hit_miss<='0';Stall<='1';
        
        when Write_Back=>
        sig_tagin<=tag;
        sig_wr<='0' ;sig_rd<='0';
      
        Cache_read<='0'; Cache_Bus_Write<='1';Memory_Bus_Read<='1';Cache_Bus_Read<='0';Memory_Bus_Write<='0';
        hit_miss<='0';Stall<='1';
        
        when Read_Main=>
        sig_tagin<=tag;
        sig_wr<='0' ;sig_rd<='0';
      
        Cache_read<='0'; Cache_Bus_Write<='0';Memory_Bus_Read<='0';Cache_Bus_Read<='1';Memory_Bus_Write<='1';
        hit_miss<='0';Stall<='1';
    end case;
end process;


end architecture ; -- arch