library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;
entity MainMemory is
  port (
    clk,rst,busRead,busWrite:IN std_logic;--bus read -->> read from bus to write to memory
    --bus write -->>  write to bus data read from memory 
    address:IN std_logic_vector(10 downto 0);
    BusDataIN:IN std_logic_vector(127 downto 0);
    BusDataOUT:OUT std_logic_vector(127 downto 0);
    counter:IN std_logic_vector(1 downto 0); -- to sync with cache.
    readySignal:Out std_logic
  ) ;
end MainMemory ;

architecture memoryARch of MainMemory is
signal WR,RD :std_logic;
signal actualAddress:std_logic_vector(10 downto 0);
signal DataIn,DataOut:std_logic_vector(31 downto 0);
begin

Actualaddress<= std_logic_vector((unsigned(counter)*2)+unsigned(address));
WR<=busRead;
RD<=busWrite;

DataIn<=BusDataIN(31 downto 0) when counter="00" and busRead ='1' else
BusDataIN(63 downto 32) when counter="01" and busRead ='1' else
BusDataIN(95 downto 64) when counter="10" and busRead ='1' else
BusDataIN(127 downto 96) when counter="11" and busRead ='1';


BusDataOUT(31 downto 0)<=DataOut  when counter="00" and busWrite='1';
BusDataOUT(63 downto 32)<=DataOut  when counter="01" and busWrite='1';
BusDataOUT(95 downto 64)<=DataOut  when counter="10" and busWrite='1';
BusDataOUT(127 downto 96)<=DataOut  when counter="11" and busWrite='1';

readySignal <= '1' when counter ="11" else '0';

MainMemory: entity work.memorymain generic map(addressBits=>11) port map (CLK=>clk,W=>WR,R=>RD,address=>Actualaddress,
dataIn=>DataIn,dataOut=>DataOut);


end architecture ; -- arch